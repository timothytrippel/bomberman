module basic_reduction(input [3:0] a, output o);
	assign o = &a;
endmodule
