module basic_constant(output [3:0] o);
	assign o = 4'b1010;
endmodule
