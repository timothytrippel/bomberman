module basic_add(input [1:0] a, input [1:0] b, output [1:0] o);
	assign o = a + b;
endmodule
