module basic_compare_eeq(input [1:0] a, input[1:0] b, output o);
	assign o = a === b;
endmodule
