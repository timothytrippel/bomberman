module constant_in_or(input b, output c);
	assign c = 1 | b;
endmodule
