module constant_in_or(input b, output c);
	assign c = b | 1;
endmodule
