module constant_part_select_pv(output [3:0] out);
	assign out[3:2] = 2'b11;
endmodule
