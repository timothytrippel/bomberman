module basic_part_select_vp(input [5:0] in, output [1:0] out);
	assign out = in[2:1];
endmodule
