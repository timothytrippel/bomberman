module padded_add(input a, input b, output [1:0] o);
	assign o = a + b;
endmodule
