module basic_part_select_pv(input [1:0] in, output [3:0] out);
	assign out[3:2] = in;
endmodule
